// ═══════════════════════════════════════════════════════════════════════════════
// NX-MIMOSA Q-TABLE WAVEFORM AGILITY MODULE
// ═══════════════════════════════════════════════════════════════════════════════
//
// Fixed-point Q-table lookup for RL-based frequency agility.
// Discretized policy from PPO agent for ultra-low latency (<10 ns @ 400 MHz).
//
// Architecture:
//   - State input: Discretized [tx_offset, jammer_estimate]
//   - Q-table: BRAM-based lookup with parallel action comparison
//   - Output: Optimal action (frequency offset) in Q8.8 format
//
// Traceability:
//   [REQ-RL-FIXED-001] Fixed-point Q-table for FPGA
//   [REQ-RL-MIT-001] Jammer mitigation via RL policy
//   [REQ-ECCM-RL] RL-based ECCM
//
// Author: Dr. Mladen Mešter / Nexellum d.o.o.
// Version: 1.1.0
// License: AGPL v3 / Commercial
// ═══════════════════════════════════════════════════════════════════════════════

`timescale 1ns/1ps

module q_table_agility #(
    // ═══════════════════════════════════════════════════════════════════════════
    // Parameters
    // ═══════════════════════════════════════════════════════════════════════════
    parameter int STATE_BITS     = 4,    // 16 discretized states per dimension
    parameter int ACTION_BITS    = 3,    // 8 discretized actions
    parameter int Q_WIDTH        = 16,   // Q8.8 signed fixed-point
    parameter int DATA_WIDTH     = 16,   // Input data width (Q8.8)
    
    // Derived parameters
    parameter int N_STATES       = (1 << STATE_BITS),
    parameter int N_ACTIONS      = (1 << ACTION_BITS),
    parameter int TABLE_SIZE     = N_STATES * N_STATES,
    
    // Action scaling (Q8.8 format)
    // Maps action index [0, N_ACTIONS-1] to freq offset [-1, +1]
    parameter logic signed [DATA_WIDTH-1:0] ACTION_MIN = -16'sd256,  // -1.0 in Q8.8
    parameter logic signed [DATA_WIDTH-1:0] ACTION_MAX = 16'sd256    // +1.0 in Q8.8
)(
    // ═══════════════════════════════════════════════════════════════════════════
    // Clock & Reset
    // ═══════════════════════════════════════════════════════════════════════════
    input  logic                          clk,
    input  logic                          rst_n,
    
    // ═══════════════════════════════════════════════════════════════════════════
    // State Input (from sensors/estimators)
    // ═══════════════════════════════════════════════════════════════════════════
    input  logic                          state_valid,
    input  logic signed [DATA_WIDTH-1:0]  state_tx_offset,      // Current TX offset (Q8.8)
    input  logic signed [DATA_WIDTH-1:0]  state_jammer_est,     // Estimated jammer freq (Q8.8)
    output logic                          state_ready,
    
    // ═══════════════════════════════════════════════════════════════════════════
    // Action Output (to waveform generator)
    // ═══════════════════════════════════════════════════════════════════════════
    output logic                          action_valid,
    output logic signed [DATA_WIDTH-1:0]  action_freq_offset,   // Optimal freq offset (Q8.8)
    output logic [ACTION_BITS-1:0]        action_index,         // Discrete action index
    input  logic                          action_ready,
    
    // ═══════════════════════════════════════════════════════════════════════════
    // Configuration & Debug
    // ═══════════════════════════════════════════════════════════════════════════
    input  logic                          cfg_enable,
    input  logic                          cfg_exploration_en,   // Enable ε-greedy exploration
    input  logic [7:0]                    cfg_epsilon,          // Exploration rate (0-255)
    input  logic [15:0]                   cfg_lfsr_seed,        // LFSR seed for randomness
    
    // Statistics
    output logic [31:0]                   stat_lookups,
    output logic [31:0]                   stat_explorations
);

    // ═══════════════════════════════════════════════════════════════════════════
    // Q-Table Memory
    // ═══════════════════════════════════════════════════════════════════════════
    // Format: q_table[state1_idx][state2_idx] = best_action_index
    // Stored as BRAM, initialized from .hex file
    
    (* ram_style = "block" *)
    logic [ACTION_BITS-1:0] q_table [0:TABLE_SIZE-1];
    
    // Initialize from file (generated by Python export)
    initial begin
        $readmemh("ppo_qtable.hex", q_table);
    end
    
    // Action value LUT (maps action index to Q8.8 offset)
    logic signed [DATA_WIDTH-1:0] action_values [0:N_ACTIONS-1];
    
    generate
        for (genvar i = 0; i < N_ACTIONS; i++) begin : gen_action_values
            // Linear interpolation: action_value = min + i * (max - min) / (N_ACTIONS - 1)
            localparam logic signed [31:0] range = ACTION_MAX - ACTION_MIN;
            localparam logic signed [31:0] scaled = ACTION_MIN + (range * i) / (N_ACTIONS - 1);
            assign action_values[i] = scaled[DATA_WIDTH-1:0];
        end
    endgenerate
    
    // ═══════════════════════════════════════════════════════════════════════════
    // LFSR for Exploration
    // ═══════════════════════════════════════════════════════════════════════════
    logic [15:0] lfsr;
    logic lfsr_bit;
    
    assign lfsr_bit = lfsr[15] ^ lfsr[14] ^ lfsr[12] ^ lfsr[3];
    
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            lfsr <= cfg_lfsr_seed;
        end else begin
            lfsr <= {lfsr[14:0], lfsr_bit};
        end
    end
    
    // ═══════════════════════════════════════════════════════════════════════════
    // Pipeline Registers
    // ═══════════════════════════════════════════════════════════════════════════
    
    // Stage 1: State discretization
    logic                          s1_valid;
    logic [STATE_BITS-1:0]         s1_state_idx_1;
    logic [STATE_BITS-1:0]         s1_state_idx_2;
    logic [$clog2(TABLE_SIZE)-1:0] s1_table_addr;
    
    // Stage 2: Table lookup
    logic                          s2_valid;
    logic [ACTION_BITS-1:0]        s2_best_action;
    logic                          s2_explore;
    
    // Stage 3: Action selection
    logic                          s3_valid;
    logic [ACTION_BITS-1:0]        s3_action_idx;
    logic signed [DATA_WIDTH-1:0]  s3_action_value;
    
    // ═══════════════════════════════════════════════════════════════════════════
    // Flow Control
    // ═══════════════════════════════════════════════════════════════════════════
    assign state_ready = cfg_enable && (!action_valid || action_ready);
    
    // ═══════════════════════════════════════════════════════════════════════════
    // STAGE 1: State Discretization
    // ═══════════════════════════════════════════════════════════════════════════
    
    function automatic logic [STATE_BITS-1:0] discretize_state(
        input logic signed [DATA_WIDTH-1:0] value
    );
        // Map Q8.8 value in [-1, +1] to [0, N_STATES-1]
        // value_normalized = (value + 256) / 512 * N_STATES
        logic signed [DATA_WIDTH+STATE_BITS:0] normalized;
        normalized = (value + 16'sd256) * N_STATES;
        return normalized[DATA_WIDTH+STATE_BITS-1:DATA_WIDTH+1];
    endfunction
    
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            s1_valid <= 1'b0;
        end else if (cfg_enable && state_valid && state_ready) begin
            s1_valid <= 1'b1;
            
            // Discretize both state components
            s1_state_idx_1 <= discretize_state(state_tx_offset);
            s1_state_idx_2 <= discretize_state(state_jammer_est);
            
            // Compute table address
            s1_table_addr <= discretize_state(state_tx_offset) * N_STATES + 
                            discretize_state(state_jammer_est);
        end else begin
            s1_valid <= 1'b0;
        end
    end
    
    // ═══════════════════════════════════════════════════════════════════════════
    // STAGE 2: Q-Table Lookup
    // ═══════════════════════════════════════════════════════════════════════════
    
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            s2_valid <= 1'b0;
            s2_explore <= 1'b0;
        end else if (s1_valid) begin
            s2_valid <= 1'b1;
            
            // BRAM lookup
            s2_best_action <= q_table[s1_table_addr];
            
            // ε-greedy exploration decision
            s2_explore <= cfg_exploration_en && (lfsr[7:0] < cfg_epsilon);
        end else begin
            s2_valid <= 1'b0;
        end
    end
    
    // ═══════════════════════════════════════════════════════════════════════════
    // STAGE 3: Action Selection
    // ═══════════════════════════════════════════════════════════════════════════
    
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            s3_valid <= 1'b0;
            s3_action_idx <= '0;
            s3_action_value <= '0;
        end else if (s2_valid) begin
            s3_valid <= 1'b1;
            
            if (s2_explore) begin
                // Random exploration: use LFSR for random action
                s3_action_idx <= lfsr[ACTION_BITS-1:0];
            end else begin
                // Exploitation: use Q-table best action
                s3_action_idx <= s2_best_action;
            end
        end else begin
            s3_valid <= 1'b0;
        end
    end
    
    // Action value lookup (combinatorial from action index)
    always_comb begin
        s3_action_value = action_values[s3_action_idx];
    end
    
    // ═══════════════════════════════════════════════════════════════════════════
    // Output Generation
    // ═══════════════════════════════════════════════════════════════════════════
    
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            action_valid <= 1'b0;
            action_freq_offset <= '0;
            action_index <= '0;
        end else if (s3_valid) begin
            action_valid <= 1'b1;
            action_freq_offset <= s3_action_value;
            action_index <= s3_action_idx;
        end else if (action_ready) begin
            action_valid <= 1'b0;
        end
    end
    
    // ═══════════════════════════════════════════════════════════════════════════
    // Statistics
    // ═══════════════════════════════════════════════════════════════════════════
    
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            stat_lookups <= '0;
            stat_explorations <= '0;
        end else begin
            if (s2_valid) begin
                stat_lookups <= stat_lookups + 1;
                if (s2_explore) begin
                    stat_explorations <= stat_explorations + 1;
                end
            end
        end
    end

endmodule


// ═══════════════════════════════════════════════════════════════════════════════
// WAVEFORM CONTROLLER WITH RL POLICY
// ═══════════════════════════════════════════════════════════════════════════════
// Top-level module integrating Q-table with DDS/NCO control

module rl_waveform_controller #(
    parameter int FREQ_WIDTH = 32,      // DDS phase accumulator width
    parameter int DATA_WIDTH = 16       // Q8.8 data width
)(
    input  logic                          clk,
    input  logic                          rst_n,
    
    // Jammer estimator interface
    input  logic                          jammer_valid,
    input  logic signed [DATA_WIDTH-1:0]  jammer_freq_est,      // Estimated jammer freq
    
    // Current waveform state
    input  logic signed [DATA_WIDTH-1:0]  current_tx_offset,
    
    // DDS/NCO control output
    output logic                          dds_update,
    output logic [FREQ_WIDTH-1:0]         dds_freq_word,
    output logic signed [DATA_WIDTH-1:0]  dds_freq_offset,
    
    // Configuration
    input  logic                          cfg_enable,
    input  logic [FREQ_WIDTH-1:0]         cfg_center_freq,      // Center frequency word
    input  logic [DATA_WIDTH-1:0]         cfg_freq_span,        // Max frequency deviation
    input  logic [15:0]                   cfg_update_interval,  // Update rate (clock cycles)
    input  logic                          cfg_exploration_en,
    input  logic [7:0]                    cfg_epsilon
);

    // ═══════════════════════════════════════════════════════════════════════════
    // Internal Signals
    // ═══════════════════════════════════════════════════════════════════════════
    
    logic                          q_action_valid;
    logic signed [DATA_WIDTH-1:0]  q_action_offset;
    logic [2:0]                    q_action_index;
    
    logic [15:0]                   update_counter;
    logic                          trigger_update;
    
    // ═══════════════════════════════════════════════════════════════════════════
    // Update Rate Control
    // ═══════════════════════════════════════════════════════════════════════════
    
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            update_counter <= '0;
            trigger_update <= 1'b0;
        end else if (cfg_enable) begin
            if (update_counter >= cfg_update_interval) begin
                update_counter <= '0;
                trigger_update <= jammer_valid;  // Only update when we have fresh jammer estimate
            end else begin
                update_counter <= update_counter + 1;
                trigger_update <= 1'b0;
            end
        end else begin
            update_counter <= '0;
            trigger_update <= 1'b0;
        end
    end
    
    // ═══════════════════════════════════════════════════════════════════════════
    // Q-Table Instance
    // ═══════════════════════════════════════════════════════════════════════════
    
    q_table_agility #(
        .STATE_BITS(4),
        .ACTION_BITS(3),
        .Q_WIDTH(16),
        .DATA_WIDTH(DATA_WIDTH)
    ) u_q_table (
        .clk(clk),
        .rst_n(rst_n),
        
        .state_valid(trigger_update),
        .state_tx_offset(current_tx_offset),
        .state_jammer_est(jammer_freq_est),
        .state_ready(),
        
        .action_valid(q_action_valid),
        .action_freq_offset(q_action_offset),
        .action_index(q_action_index),
        .action_ready(1'b1),
        
        .cfg_enable(cfg_enable),
        .cfg_exploration_en(cfg_exploration_en),
        .cfg_epsilon(cfg_epsilon),
        .cfg_lfsr_seed(16'hACE1),
        
        .stat_lookups(),
        .stat_explorations()
    );
    
    // ═══════════════════════════════════════════════════════════════════════════
    // DDS Control
    // ═══════════════════════════════════════════════════════════════════════════
    
    logic signed [FREQ_WIDTH-1:0] freq_offset_scaled;
    
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            dds_update <= 1'b0;
            dds_freq_word <= '0;
            dds_freq_offset <= '0;
        end else if (q_action_valid) begin
            // Scale Q8.8 offset to frequency word
            // offset_scaled = action_offset * freq_span / 256
            freq_offset_scaled = (q_action_offset * $signed({1'b0, cfg_freq_span})) >>> 8;
            
            dds_freq_word <= cfg_center_freq + freq_offset_scaled;
            dds_freq_offset <= q_action_offset;
            dds_update <= 1'b1;
        end else begin
            dds_update <= 1'b0;
        end
    end

endmodule


// ═══════════════════════════════════════════════════════════════════════════════
// JAMMER ESTIMATOR
// ═══════════════════════════════════════════════════════════════════════════════
// Estimates jammer frequency from power spectrum

module jammer_frequency_estimator #(
    parameter int FFT_SIZE = 1024,
    parameter int DATA_WIDTH = 16
)(
    input  logic                          clk,
    input  logic                          rst_n,
    
    // FFT magnitude input
    input  logic                          fft_valid,
    input  logic [DATA_WIDTH-1:0]         fft_magnitude,
    input  logic [$clog2(FFT_SIZE)-1:0]   fft_bin,
    input  logic                          fft_last,
    
    // Jammer estimate output
    output logic                          jammer_valid,
    output logic signed [DATA_WIDTH-1:0]  jammer_freq_est,     // Normalized [-1, +1]
    output logic [DATA_WIDTH-1:0]         jammer_power,        // Peak power
    output logic                          jammer_detected,
    
    // Configuration
    input  logic [DATA_WIDTH-1:0]         cfg_detection_thresh, // dB threshold
    input  logic [DATA_WIDTH-1:0]         cfg_noise_floor
);

    // Peak tracking
    logic [DATA_WIDTH-1:0]         peak_power;
    logic [$clog2(FFT_SIZE)-1:0]   peak_bin;
    logic [DATA_WIDTH-1:0]         power_sum;
    logic [$clog2(FFT_SIZE)-1:0]   bin_count;
    
    // Processing
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            peak_power <= '0;
            peak_bin <= '0;
            power_sum <= '0;
            bin_count <= '0;
            jammer_valid <= 1'b0;
            jammer_detected <= 1'b0;
        end else if (fft_valid) begin
            // Track peak
            if (fft_magnitude > peak_power) begin
                peak_power <= fft_magnitude;
                peak_bin <= fft_bin;
            end
            
            // Accumulate for average
            power_sum <= power_sum + fft_magnitude;
            bin_count <= bin_count + 1;
            
            if (fft_last) begin
                // Output result
                jammer_valid <= 1'b1;
                jammer_power <= peak_power;
                
                // Convert bin to normalized frequency [-1, +1]
                // freq = (bin - FFT_SIZE/2) / (FFT_SIZE/2)
                jammer_freq_est <= ((peak_bin - FFT_SIZE/2) <<< 9) / (FFT_SIZE/2);
                
                // Detection: peak > threshold above noise
                jammer_detected <= (peak_power > cfg_noise_floor + cfg_detection_thresh);
                
                // Reset for next frame
                peak_power <= '0;
                power_sum <= '0;
                bin_count <= '0;
            end
        end else begin
            jammer_valid <= 1'b0;
        end
    end

endmodule
